library verilog;
use verilog.vl_types.all;
entity ffjk_vlg_vec_tst is
end ffjk_vlg_vec_tst;
