library verilog;
use verilog.vl_types.all;
entity fft_vlg_vec_tst is
end fft_vlg_vec_tst;
