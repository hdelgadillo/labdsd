library verilog;
use verilog.vl_types.all;
entity contador3bits_vlg_vec_tst is
end contador3bits_vlg_vec_tst;
