library verilog;
use verilog.vl_types.all;
entity contador3bits_vlg_check_tst is
    port(
        salcuenta       : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end contador3bits_vlg_check_tst;
