library verilog;
use verilog.vl_types.all;
entity miflip_vlg_vec_tst is
end miflip_vlg_vec_tst;
